module simpleand(f,x,y);
      input x,y;
      output f;
      and G1(f,x,y);
endmodule
